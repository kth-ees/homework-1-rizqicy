module csa_8 (
  input logic [7:0] a, b,
  output logic [7:0] sum,
  output logic carry
);
  // 8-bit adder with Carry Select Adder
  logic c_sel, cout0, cout1;
  logic [3:0]sum3_0;
  logic [3:0]sum_c0;
  logic [3:0]sum_c1;

  adder_4 adder0_3 (.A(a[3:0]), .B(b[3:0]), .sum(sum3_0), .carry(c_sel));
  adder_4 adder4_7_c0 (.A(a[7:4]), .B(b[7:4]), .sum(sum_c0), .carry(cout0));
  adder_4 adder4_7_c1 (.A(a[7:4]), .B((b[7:4] + 1)), .sum(sum_c1), .carry(cout1));

  assign carry = (c_sel) ? cout1 : cout0;
  assign sum = (c_sel) ? {sum_c1,sum3_0} : {sum_c0,sum3_0};

endmodule
